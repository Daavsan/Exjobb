** Profile: "SCHEMATIC1-Trans"  [ C:\Users\A1201-admin\Documents\Exjobb\Orcad\Filter Test-PSpiceFiles\SCHEMATIC1\Trans.sim ] 

** Creating circuit file "Trans.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\A1201-admin\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "C:\Users\A1201-admin\Documents\Exjobb\Orcad\lmg1210.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
