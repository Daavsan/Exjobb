** Profile: "SCHEMATIC1-trans"  [ C:\Users\A1201-admin\Documents\Exjobb\Orcad\filter-pspicefiles\schematic1\trans.sim ] 

** Creating circuit file "trans.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\A1201-admin\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "C:\Users\A1201-admin\Documents\Exjobb\Orcad\lmg1210.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 7u 0 0.1n 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
