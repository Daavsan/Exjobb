** Profile: "SCHEMATIC1-trans_1"  [ c:\users\a1201-admin\documents\exjobb\orcad\mostest_cadence-PSpiceFiles\SCHEMATIC1\trans_1.sim ] 

** Creating circuit file "trans_1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\A1201-admin\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "C:\Users\A1201-admin\Documents\Exjobb\Orcad\lmg1210.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10ns 0 
.OPTIONS ADVCONV
.AUTOCONVERGE ITL1=1000 ITL2=1000 ITL4=1000 RELTOL=0.05 ABSTOL=1.0E-6 VNTOL=.001 PIVTOL=1.0E-10 
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
